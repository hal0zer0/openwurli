* Wurlitzer 200A Preamp THD Comparison: Real Q2N5089 vs Ideal BJT
* ================================================================
* Purpose: Measure harmonic distortion at 262 Hz (C4) across 4 input
*          amplitudes, comparing the full Gummel-Poon Q2N5089 model
*          against the beta-infinity ideal model used in the DK DSP code.
*
* Circuit: Full 200A preamp with C20, D1, Rload. R_ldr = 1M (no tremolo).
*          Two identical instances: suffix _r (real) and _i (ideal).
*
* Input levels (peak amplitude at source, before R1=22K):
*   1 mV   — pp/quiet
*   10 mV  — mf/moderate
*   50 mV  — f/loud
*   100 mV — ff/clipping territory
*
* Analysis: transient 500ms, fourier from last ~78 cycles (262 Hz).
*           ngspice fourier command reports H1-H9 and THD automatically.
*
* Run: ngspice -b tb_real_thd.cir  (or ngspice -r ... for rawfile)

.title THD Comparison: Real Q2N5089 vs Ideal BJT at 262 Hz

* ==================================================================
* TRANSISTOR MODELS
* ==================================================================

* Ideal model: very high BF, no parasitics (matches DK DSP assumptions)
.MODEL Q_IDEAL NPN(
+  IS=3.03E-14 BF=100000 NF=1.0 VAF=1000
+  RB=0 RE=0 RC=0
+  CJE=0 CJC=0 TF=0 TR=0)

* Full Gummel-Poon model for 2N5089 (Fairchild)
.MODEL Q2N5089 NPN(
+  IS=3.03E-14 BF=1434 NF=1.005 VAF=98.5 IKF=0.01358
+  ISE=2.88E-15 NE=1.262 BR=4.62 NR=1 VAR=22 IKR=0.1
+  ISC=1.065E-11 NC=1.41 RB=57 RE=0.518 RC=2.58
+  CJE=3.22E-12 VJE=0.65 MJE=0.33 TF=5.4E-10
+  CJC=1.35E-12 VJC=0.4 MJC=0.33 XCJC=0.63 TR=5E-08
+  XTB=1.38 EG=1.11 XTI=3 FC=0.5)

* Diode for bias protection (real circuit only)
.MODEL D1N4148 D(IS=2.52E-09 RS=0.568 N=1.752 BV=100 IBV=100E-06
+  CJO=4E-12 VJ=0.7 M=0.45 TT=6E-09)

* ==================================================================
* CIRCUIT R: REAL Q2N5089 (full SPICE model + C20, D1, Rload)
* ==================================================================
Vcc_r   vcc_r   0   DC 15
Vin_r   src_r   0   DC 0 SIN(0 0.001 262 0 0)

* Input network
R1_r    src_r   nodeA_r   22K
Cin_r   nodeA_r base1_r   0.022U

* Bias network with C20 and D1
R2_r    vcc_r   base1_r   2MEG
R3_r    base1_r 0         470K
C20_r   base1_r 0         220P
D1_r    0       base1_r   D1N4148

* Stage 1: TR-1
Q1_r    coll1_r base1_r emit1_r Q2N5089
Rc1_r   vcc_r   coll1_r   150K
Cc3_r   coll1_r base1_r   100P
Re1_r   emit1_r 0         33K
Ce1_r   emit1_r fb_j_r    4.7U

* Feedback network (no tremolo: Rldr = 1M)
R10_r   out_r   fb_j_r    56K
Rldr_r  fb_j_r  0         1MEG

* Stage 2: TR-2
Q2_r    coll2_r coll1_r emit2a_r Q2N5089
Rc2_r   vcc_r   coll2_r   1.8K
Re2a_r  emit2a_r emit2b_r 270
Ce2_r   emit2a_r emit2b_r 22U
Re2b_r  emit2b_r 0        820
Cc4_r   coll2_r  coll1_r  100P

* Output
R9_r    coll2_r out_r     6.8K
Rload_r out_r   0         100K

* ==================================================================
* CIRCUIT I: IDEAL BJT (beta=100000, no parasitics, no C20/D1/Rload)
* ==================================================================
* Note: Keeping C20, D1, and Rload here too for apples-to-apples
* circuit topology comparison. The ONLY difference is the BJT model.
Vcc_i   vcc_i   0   DC 15
Vin_i   src_i   0   DC 0 SIN(0 0.001 262 0 0)

* Input network
R1_i    src_i   nodeA_i   22K
Cin_i   nodeA_i base1_i   0.022U

* Bias network with C20 and D1 (same topology as real)
R2_i    vcc_i   base1_i   2MEG
R3_i    base1_i 0         470K
C20_i   base1_i 0         220P
D1_i    0       base1_i   D1N4148

* Stage 1: TR-1
Q1_i    coll1_i base1_i emit1_i Q_IDEAL
Rc1_i   vcc_i   coll1_i   150K
Cc3_i   coll1_i base1_i   100P
Re1_i   emit1_i 0         33K
Ce1_i   emit1_i fb_j_i    4.7U

* Feedback network (no tremolo: Rldr = 1M)
R10_i   out_i   fb_j_i    56K
Rldr_i  fb_j_i  0         1MEG

* Stage 2: TR-2
Q2_i    coll2_i coll1_i emit2a_i Q_IDEAL
Rc2_i   vcc_i   coll2_i   1.8K
Re2a_i  emit2a_i emit2b_i 270
Ce2_i   emit2a_i emit2b_i 22U
Re2b_i  emit2b_i 0        820
Cc4_i   coll2_i  coll1_i  100P

* Output
R9_i    coll2_i out_i     6.8K
Rload_i out_i   0         100K

* ==================================================================
* SIMULATION CONTROL
* ==================================================================
.control

set filetype = ascii

echo ""
echo "================================================================="
echo "  THD COMPARISON: Real Q2N5089 vs Ideal BJT"
echo "  Frequency: 262 Hz (C4)"
echo "  Preamp: Rldr = 1M (no tremolo, gain ~2.0x)"
echo "================================================================="
echo ""

* First: verify DC operating points
op

echo "=== DC OPERATING POINT: Real Q2N5089 ==="
echo "TR-1 (expected: B=2.45V, E=1.95V, C=4.1V):"
print v(base1_r) v(emit1_r) v(coll1_r)
echo "TR-2 (expected: B=4.1V, E=3.4V, C=8.8V):"
print v(coll1_r) v(emit2a_r) v(coll2_r)
echo "Output and feedback junction:"
print v(out_r) v(fb_j_r)
echo ""

echo "=== DC OPERATING POINT: Ideal BJT ==="
echo "TR-1 (expected: B=2.45V, E=1.95V, C=4.1V):"
print v(base1_i) v(emit1_i) v(coll1_i)
echo "TR-2 (expected: B=4.1V, E=3.4V, C=8.8V):"
print v(coll1_i) v(emit2a_i) v(coll2_i)
echo "Output and feedback junction:"
print v(out_i) v(fb_j_i)
echo ""

* Reset for transient
reset

echo "================================================================="
echo "  SWEEPING INPUT AMPLITUDES"
echo "================================================================="
echo ""

* Sweep 4 amplitude levels
foreach amp_val 0.001 0.010 0.050 0.100

  * Set both sources to same amplitude
  alter @vin_r[sin] = [ 0 $amp_val 262 0 0 ]
  alter @vin_i[sin] = [ 0 $amp_val 262 0 0 ]

  * Transient: 500ms total, skip first 200ms for steady state.
  * Timestep 1us -> 262 Hz needs ~3817 us/cycle, so ~1 us gives
  * ~3817 points/cycle, more than adequate for Fourier up to H9.
  tran 1u 500m 200m 1u

  echo ""
  echo "============================================================"
  echo "  Input amplitude: $amp_val V peak at 262 Hz"
  echo "============================================================"
  echo ""

  * Output peak-to-peak measurements
  echo "--- REAL Q2N5089 ---"
  meas tran real_out_pp PP v(out_r) from=300m to=500m
  meas tran real_out_max MAX v(out_r) from=300m to=500m
  meas tran real_out_min MIN v(out_r) from=300m to=500m
  meas tran real_c1_pp PP v(coll1_r) from=300m to=500m

  echo ""
  echo "Fourier analysis — REAL preamp output:"
  fourier 262 v(out_r)

  echo ""
  echo "Fourier analysis — REAL Stage 1 collector:"
  fourier 262 v(coll1_r)

  echo ""
  echo "--- IDEAL BJT ---"
  meas tran ideal_out_pp PP v(out_i) from=300m to=500m
  meas tran ideal_out_max MAX v(out_i) from=300m to=500m
  meas tran ideal_out_min MIN v(out_i) from=300m to=500m
  meas tran ideal_c1_pp PP v(coll1_i) from=300m to=500m

  echo ""
  echo "Fourier analysis — IDEAL preamp output:"
  fourier 262 v(out_i)

  echo ""
  echo "Fourier analysis — IDEAL Stage 1 collector:"
  fourier 262 v(coll1_i)

  * Reset state for next iteration (important: keeps models intact)
  reset

end

echo ""
echo "================================================================="
echo "  ALL AMPLITUDES COMPLETE"
echo "================================================================="
echo ""

* Bonus: tremolo bright (Rldr=19K) at 50 mV to see if gain boost
* pushes the real circuit further into nonlinearity
echo ""
echo "================================================================="
echo "  BONUS: Tremolo Bright (Rldr=19K) at 50 mV peak"
echo "  Gain ~4x, so 50 mV input -> ~200 mV pp swing (vs ~100 mV no trem)"
echo "================================================================="
echo ""

* Change LDR to 19K for both circuits
alter rldr_r = 19000
alter rldr_i = 19000
alter @vin_r[sin] = [ 0 0.050 262 0 0 ]
alter @vin_i[sin] = [ 0 0.050 262 0 0 ]

tran 1u 500m 200m 1u

echo "--- REAL Q2N5089, Rldr=19K, 50mV peak ---"
meas tran real_out_pp PP v(out_r) from=300m to=500m
echo "Fourier — REAL preamp output (tremolo bright):"
fourier 262 v(out_r)

echo ""
echo "--- IDEAL BJT, Rldr=19K, 50mV peak ---"
meas tran ideal_out_pp PP v(out_i) from=300m to=500m
echo "Fourier — IDEAL preamp output (tremolo bright):"
fourier 262 v(out_i)

echo ""
echo "================================================================="
echo "  TESTBENCH COMPLETE"
echo "================================================================="

quit

.endc
.end
