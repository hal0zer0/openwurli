.title Wurlitzer 200A Preamp - Topology B LDR Sweep
* Test emitter feedback topology with correct LDR path resistances
* LDR path includes: 18K + 680 + LDR_resistance
* So minimum path resistance ~19K (LDR fully bright)
* Maximum path resistance ~1MEG (LDR fully dark / tremolo off)

.MODEL Q2N5089 NPN(
+  IS=3.03E-14 BF=1434 NF=1.005 VAF=98.5 IKF=0.01358
+  ISE=2.88E-15 NE=1.262 BR=4.62 NR=1 VAR=22 IKR=0.1
+  ISC=1.065E-11 NC=1.41 RB=57 RE=0.518 RC=2.58
+  CJE=3.22E-12 VJE=0.65 MJE=0.33 TF=5.4E-10
+  CJC=1.35E-12 VJC=0.4 MJC=0.33 XCJC=0.63 TR=5E-08
+  XTB=1.38 EG=1.11 XTI=3 FC=0.5)
.MODEL D1N4148 D(IS=2.52E-09 RS=0.568 N=1.752 BV=100
+  IBV=100E-06 CJO=4E-12 VJ=0.7 M=0.45 TT=6E-09)

Vcc vcc 0 DC 15

* Preamp with emitter feedback topology
Vin in_sig 0 DC 0 SIN(0 0.002 440)
R1 in_sig node_A 22K
Cin node_A base1 0.022U
R2 vcc base1 2MEG
R3 base1 0 470K
C20 base1 0 220P
D1 0 base1 D1N4148
Q1 coll1 base1 emit1 Q2N5089
Rc1 vcc coll1 150K
Cc3 coll1 base1 100P
Re1 emit1 0 33K
Ce1 emit1 fb_junct 4.7U
Q2 coll2 coll1 emit2a Q2N5089
Rc2 vcc coll2 1.8K
Re2a emit2a emit2b 270
Ce2 emit2a emit2b 22U
Re2b emit2b 0 820
Cc4 coll2 coll1 100P
R9 coll2 out 6.8K
Rload out 0 100K
R10 out fb_junct 56K
Rldr_path fb_junct 0 19K

.control
echo "============================================================"
echo "TOPOLOGY B: LDR SWEEP (emitter feedback)"
echo "Input: 2mV peak at 440 Hz"
echo "============================================================"
echo ""

* Sweep LDR path resistance from 19K (full bright) to 1MEG (off)
* Values chosen to span realistic tremolo range

foreach rldr_val 19K 25K 33K 47K 68K 100K 150K 220K 330K 470K 680K 1MEG
  alter Rldr_path = $rldr_val
  destroy all
  tran 0.5u 200m
  meas tran vmax max v(out) from=150m to=200m
  meas tran vmin min v(out) from=150m to=200m
  meas tran vc1max max v(coll1) from=150m to=200m
  meas tran vc1min min v(coll1) from=150m to=200m
  fourier 440 v(out)
  echo ""
end

echo "============================================================"
echo "ADDITIONAL: Test different input levels at key Rldr values"
echo "============================================================"

* --- 19K (tremolo bright), mf level ---
echo ""
echo "=== Rldr=19K (bright), various inputs ==="
alter Rldr_path = 19K

foreach amp_val 0.0005 0.001 0.002 0.005 0.010 0.050
  alter Vin DC=0 AC=0 SIN 0 $amp_val 440
  destroy all
  tran 0.5u 200m
  meas tran vmax max v(out) from=150m to=200m
  meas tran vmin min v(out) from=150m to=200m
  fourier 440 v(out)
  echo ""
end

* --- 1MEG (no tremolo), various inputs ---
echo ""
echo "=== Rldr=1MEG (dark/off), various inputs ==="
alter Rldr_path = 1MEG

foreach amp_val 0.0005 0.001 0.002 0.005 0.010 0.050
  alter Vin DC=0 AC=0 SIN 0 $amp_val 440
  destroy all
  tran 0.5u 200m
  meas tran vmax max v(out) from=150m to=200m
  meas tran vmin min v(out) from=150m to=200m
  fourier 440 v(out)
  echo ""
end

echo "============================================================"
echo "SWEEP COMPLETE"
echo "============================================================"

.endc
.end
