* Wurlitzer 200A Preamp — Tremolo Pump DC Analysis
* ================================================
* Measures:
*   1. DC operating point at V(out) as R_ldr varies from 1M to 19K
*   2. Transient response showing the multi-volt DC swing during tremolo
*   3. What C-8 (4.7uF) into R-31 (15K) does to the pump signal
*
* This testbench answers: "Is the multi-volt DC swing at V(out) real physics,
* or a modeling artifact?"

.title Preamp Pump Analysis - DC Sweep and Transient

.include ../models/transistors.lib
.include ../models/diodes.lib
.include ../subcircuits/preamp.cir

* Supply
Vcc  vcc 0  DC 15

* Instantiate preamp
Xpre  in_sig out vcc 0 fb_junct  wurli_preamp

* No audio signal -- just measure pump from R_ldr modulation
R1   in_sig 0  22K
* R-1 in the real circuit goes to the pickup plate (150V through 1M feed);
* for pump analysis we ground it through R1 to isolate the pump source.

* === Test 1: DC Sweep of R_ldr ===
* Sweep a resistor from fb_junct to ground.
* We use a voltage source + resistor to parametrize.
* Actually, for DC sweep we just do multiple .OP runs via parameter.

* For DC operating point analysis, use a fixed R_ldr:
* R_ldr_path = 19K (tremolo bright peak)
Rldr_bright  fb_junct 0  19K

.OP

.end
