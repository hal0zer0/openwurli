.title Wurlitzer 200A Preamp - AC Sweep (Corrected Emitter Feedback)
* Measures closed-loop gain and bandwidth with corrected topology
* R-10 feeds back from output to TR-1 emitter via Ce1 (4.7uF coupling cap)

.MODEL Q2N5089 NPN(
+  IS=3.03E-14 BF=1434 NF=1.005 VAF=98.5 IKF=0.01358
+  ISE=2.88E-15 NE=1.262 BR=4.62 NR=1 VAR=22 IKR=0.1
+  ISC=1.065E-11 NC=1.41 RB=57 RE=0.518 RC=2.58
+  CJE=3.22E-12 VJE=0.65 MJE=0.33 TF=5.4E-10
+  CJC=1.35E-12 VJC=0.4 MJC=0.33 XCJC=0.63 TR=5E-08
+  XTB=1.38 EG=1.11 XTI=3 FC=0.5)

.MODEL D1N4148 D(IS=2.52E-09 RS=0.568 N=1.752 BV=100
+  IBV=100E-06 CJO=4E-12 VJ=0.7 M=0.45 TT=6E-09)

Vcc vcc 0 DC 15

* Input signal source through R1 (22K) - represents reed bar pickup
Vin in_sig 0 DC 0 AC 1
R1 in_sig node_A 22K

* Input coupling to base1
Cin node_A base1 0.022U

* Base1 bias and filtering
R2 vcc base1 2MEG
R3 base1 0 470K
C20 base1 0 220P
D1 0 base1 D1N4148

* Stage 1: TR-1
Q1 coll1 base1 emit1 Q2N5089
Rc1 vcc coll1 150K
Cc3 coll1 base1 100P

* TR-1 emitter: Re1 to ground (DC path), Ce1 to feedback junction (AC coupling)
Re1 emit1 0 33K
Ce1 emit1 fb_junct 4.7U

* Feedback junction: R-10 from output, Ce1 to emitter, LDR path to ground
* Rldr_path = 50K vibrato (assume mid position ~25K) + 18K + LDR_dark (~100K+)
* For no-tremolo baseline: LDR is dark, very high resistance
* Model as 120K total (conservative estimate for LDR dark path)
Rldr_path fb_junct 0 120K

* R-10 feedback from output to junction
R10 out fb_junct 56K

* Stage 2: TR-2 (direct-coupled from coll1)
Q2 coll2 coll1 emit2a Q2N5089
Rc2 vcc coll2 1.8K
Re2a emit2a emit2b 270
Ce2 emit2a emit2b 22U
Re2b emit2b 0 820
Cc4 coll2 coll1 100P

* Output
R9 coll2 out 6.8K
Rload out 0 100K

.control
* DC operating point first
op
echo "=== DC Operating Point ==="
print v(base1) v(emit1) v(coll1) v(coll2) v(fb_junct) v(out)
print @q1[ic] @q2[ic] @q1[gm] @q2[gm]

* AC sweep: 1 Hz to 1 MHz, 200 points per decade
ac dec 200 1 1MEG

* Write full frequency response data
* Vin = 1V AC, so vdb(out) IS the gain in dB directly
wrdata /tmp/preamp_ac_gain.txt vdb(out) vp(out) vdb(base1) vdb(emit1) vdb(fb_junct) vdb(coll1) vdb(coll2)

* Find and print key measurements
echo ""
echo "=== Gain at Key Frequencies ==="
echo "Format: frequency, gain_dB, gain_linear"
let gain_db = vdb(out)
let gain_lin = vm(out)

* Print gain at specific frequencies
print gain_db[200] gain_lin[200]
* ~100 Hz (index varies - use meas)
meas ac gain_100 find vdb(out) at=100
meas ac gain_1k find vdb(out) at=1000
meas ac gain_2k find vdb(out) at=2000
meas ac gain_5k find vdb(out) at=5000
meas ac gain_10k find vdb(out) at=10000
meas ac gain_20k find vdb(out) at=20000

* Find peak gain
meas ac peak_gain max vdb(out)
meas ac peak_freq max_at vdb(out)

* Find -3dB bandwidth (relative to peak)
let target = peak_gain - 3
meas ac bw_low when vdb(out)=target rise=1
meas ac bw_high when vdb(out)=target fall=last

echo ""
echo "=== Summary ==="

.endc

.end
