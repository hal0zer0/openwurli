.title Wurlitzer 200A Preamp - Corrected Emitter Feedback Topology
* R-10 feeds back from output to TR-1 emitter via Ce1 (4.7uF coupling cap)
* Re1 (33K) provides separate DC path from emitter to ground
* Ce1 AC-couples the feedback junction to the emitter
* This is NEGATIVE feedback (series-series / emitter feedback)

.MODEL Q2N5089 NPN(
+  IS=3.03E-14 BF=1434 NF=1.005 VAF=98.5 IKF=0.01358
+  ISE=2.88E-15 NE=1.262 BR=4.62 NR=1 VAR=22 IKR=0.1
+  ISC=1.065E-11 NC=1.41 RB=57 RE=0.518 RC=2.58
+  CJE=3.22E-12 VJE=0.65 MJE=0.33 TF=5.4E-10
+  CJC=1.35E-12 VJC=0.4 MJC=0.33 XCJC=0.63 TR=5E-08
+  XTB=1.38 EG=1.11 XTI=3 FC=0.5)

.MODEL D1N4148 D(IS=2.52E-09 RS=0.568 N=1.752 BV=100
+  IBV=100E-06 CJO=4E-12 VJ=0.7 M=0.45 TT=6E-09)

Vcc vcc 0 DC 15

* Input signal source through R1 (22K) - represents reed bar pickup
Vin in_sig 0 DC 0 AC 0.01
R1 in_sig node_A 22K

* Input coupling to base1
Cin node_A base1 0.022U

* Base1 bias and filtering
R2 vcc base1 2MEG
R3 base1 0 470K
C20 base1 0 220P
D1 0 base1 D1N4148

* Stage 1: TR-1
Q1 coll1 base1 emit1 Q2N5089
Rc1 vcc coll1 150K
Cc3 coll1 base1 100P

* TR-1 emitter: Re1 to ground (DC path), Ce1 to feedback junction (AC coupling)
Re1 emit1 0 33K
Ce1 emit1 fb_junct 4.7U

* Feedback junction: R-10 from output, Ce1 to emitter, ground path
* In real circuit, DC ground for this node is through Pin 1 -> cable -> LDR -> ground
* For now, model with a large resistor to ground (LDR dark = high resistance)
* LDR path: 18K + 680 + LDR (model as Rldr variable)
Rldr_path fb_junct 0 120K

* R-10 feedback from output to junction
R10 out fb_junct 56K

* Stage 2: TR-2 (direct-coupled from coll1)
Q2 coll2 coll1 emit2a Q2N5089
Rc2 vcc coll2 1.8K
Re2a emit2a emit2b 270
Ce2 emit2a emit2b 22U
Re2b emit2b 0 820
Cc4 coll2 coll1 100P

* Output
R9 coll2 out 6.8K
Rload out 0 100K

.control
* DC operating point
op
print v(node_A) v(base1) v(emit1) v(fb_junct) v(coll1) v(coll2) v(out)

* Transient - check for stability (no input signal)
tran 10u 50m
wrdata /tmp/emitter_fb_tran.txt v(node_A) v(base1) v(emit1) v(fb_junct) v(coll1) v(coll2) v(out)

* AC sweep
ac dec 100 10 100K
wrdata /tmp/emitter_fb_ac.txt vdb(out) vp(out) vdb(base1) vdb(emit1) vdb(fb_junct)
.endc

.end
