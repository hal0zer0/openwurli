* Wurlitzer 200A Preamp — DC Operating Point vs R_ldr (compact output)
* ===================================================================

.title Preamp DC vs R_ldr - Compact

.include ../models/transistors.lib
.include ../models/diodes.lib
.include ../subcircuits/preamp.cir

* Supply
Vcc  vcc 0  DC 15

* Instantiate preamp
Xpre  in_sig out vcc 0 fb_junct  wurli_preamp

* No audio — ground input
Vin  in_sig 0  DC 0

* LDR path: parametric sweep
Vldr_ctrl  ldr_ctrl 0  DC 19K
Rldr  fb_junct 0  R='V(ldr_ctrl)'

* Sweep R_ldr from 19K to 1M in larger steps for readable output
.DC Vldr_ctrl 19K 1000K 100K

* Only print the key nodes
.print DC V(out) V(fb_junct)

.end
